module constants

// PVNO is the Protocol Version Number.
// See https://datatracker.ietf.org/doc/html/rfc4120#section-7.5.6
pub const pvno = 5
