module vkerberos

const vkerberos_version = '0.1.0'