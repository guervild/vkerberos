module types

// https://datatracker.ietf.org/doc/html/rfc4120#section-5.2.6
// pub struct AuthorizationDataEntry {
// pub mut:
// 	ad_type int
// 	ad_data []u8
// }

// type AuthorizationData = []AuthorizationDataEntry

// type ADIfRelevant = AuthorizationData
