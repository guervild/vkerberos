module types

pub const kdcflagsreserved = int(0)
pub const kdcflagsforwardable = int(1)
pub const kdcflagsforwarded = int(2)
pub const kdcflagsproxiable = int(3)
pub const kdcflagsproxy = int(4)
pub const kdcflagsallowpostdate = int(5)
pub const kdcflagspostdated = int(6)
pub const kdcflagsrenewable = int(8)
pub const kdcflagsopthardwareauth = int(11)
pub const kdcflagsconstraineddelegation = int(14)
pub const kdcflagscanonicalize = int(15)
pub const kdcflagsrequestanonymous = int(16)
pub const kdcflagscnameinadditionalticket = int(17)
pub const kdcflagsdisabletransitedcheck = int(26)
pub const kdcflagsrenewableok = int(27)
pub const kdcflagsenctktinskey = int(28)
pub const kdcflagsrenew = int(30)
pub const kdcflagsvalidate = int(31)
